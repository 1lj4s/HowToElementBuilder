* EQUIVALENT CIRCUIT FOR VECTOR FITTED S-MATRIX
* Created using scikit-rf vectorFitting.py
*
.SUBCKT s_equivalent p1 p2
*
* Port network for port 1
V1 p1 s1 0
R1 s1 0 50.0
Gd1_1 0 s1 p1 0 -0.05599437861010731
Fd1_1 0 s1 V1 -2.7997189305053656
Gr1_1_1 0 s1 x1_a1 0 3749671826091.7427
Gr2_re_1_1 0 s1 x2_re_a1 0 -20119730888.36101
Gr2_im_1_1 0 s1 x2_im_a1 0 -7615793267.56339
Gr3_re_1_1 0 s1 x3_re_a1 0 -4582270774.515794
Gr3_im_1_1 0 s1 x3_im_a1 0 327605610.7607881
Gr4_re_1_1 0 s1 x4_re_a1 0 -4687608450.879957
Gr4_im_1_1 0 s1 x4_im_a1 0 -60815242.74458452
Gr5_re_1_1 0 s1 x5_re_a1 0 -4703207822.656034
Gr5_im_1_1 0 s1 x5_im_a1 0 -73675770.72488609
Gr6_re_1_1 0 s1 x6_re_a1 0 -4696210203.28238
Gr6_im_1_1 0 s1 x6_im_a1 0 -70184505.16911012
Gr7_re_1_1 0 s1 x7_re_a1 0 -4690028374.353796
Gr7_im_1_1 0 s1 x7_im_a1 0 -82816399.82581234
Gr8_re_1_1 0 s1 x8_re_a1 0 -4721421341.403379
Gr8_im_1_1 0 s1 x8_im_a1 0 -106419878.93335082
Gr9_1_1 0 s1 x9_a1 0 -4689776981.4304285
Gr10_re_1_1 0 s1 x10_re_a1 0 1043910.4473995286
Gr10_im_1_1 0 s1 x10_im_a1 0 -118841.77270054491
Gr11_1_1 0 s1 x11_a1 0 4592739.71891656
Gd1_2 0 s1 p2 0 -0.0016856930057704883
Fd1_2 0 s1 V2 -0.08428465028852442
Gr1_1_2 0 s1 x1_a2 0 114980691786.52382
Gr2_re_1_2 0 s1 x2_re_a2 0 -3439807808.4147644
Gr2_im_1_2 0 s1 x2_im_a2 0 2514561760.7023377
Gr3_re_1_2 0 s1 x3_re_a2 0 4423321369.53323
Gr3_im_1_2 0 s1 x3_im_a2 0 -651374200.6221427
Gr4_re_1_2 0 s1 x4_re_a2 0 -4684893909.527276
Gr4_im_1_2 0 s1 x4_im_a2 0 -61217124.35522651
Gr5_re_1_2 0 s1 x5_re_a2 0 4712777508.873276
Gr5_im_1_2 0 s1 x5_im_a2 0 73744102.59193671
Gr6_re_1_2 0 s1 x6_re_a2 0 -4702204173.996921
Gr6_im_1_2 0 s1 x6_im_a2 0 -68486113.03858867
Gr7_re_1_2 0 s1 x7_re_a2 0 4691734541.675555
Gr7_im_1_2 0 s1 x7_im_a2 0 92677089.01510376
Gr8_re_1_2 0 s1 x8_re_a2 0 -4725312491.31795
Gr8_im_1_2 0 s1 x8_im_a2 0 -120007193.34835783
Gr9_1_2 0 s1 x9_a2 0 4665975028.099103
Gr10_re_1_2 0 s1 x10_re_a2 0 -560743.618316202
Gr10_im_1_2 0 s1 x10_im_a2 0 2135652.8297406496
Gr11_1_2 0 s1 x11_a2 0 -1099763.15568693
*
* State networks driven by port 1
Cx1_a1 x1_a1 0 1.0
Gx1_a1 0 x1_a1 p1 0 0.07071067811865475
Fx1_a1 0 x1_a1 V1 3.5355339059327378
Rp1_a1 0 x1_a1 3.1658774695127977e-13
Cx2_re_a1 x2_re_a1 0 1.0
Gx2_re_a1 0 x2_re_a1 p1 0 0.1414213562373095
Fx2_re_a1 0 x2_re_a1 V1 7.0710678118654755
Rp2_re_re_a1 0 x2_re_a1 3.094780737837525e-11
Gp2_re_im_a1 0 x2_re_a1 x2_im_a1 0 338816889165.91437
Cx2_im_a1 x2_im_a1 0 1.0
Gp2_im_re_a1 0 x2_im_a1 x2_re_a1 0 -338816889165.91437
Rp2_im_im_a1 0 x2_im_a1 3.094780737837525e-11
Cx3_re_a1 x3_re_a1 0 1.0
Gx3_re_a1 0 x3_re_a1 p1 0 0.1414213562373095
Fx3_re_a1 0 x3_re_a1 V1 7.0710678118654755
Rp3_re_re_a1 0 x3_re_a1 6.71721917054064e-11
Gp3_re_im_a1 0 x3_re_a1 x3_im_a1 0 262327540913.7152
Cx3_im_a1 x3_im_a1 0 1.0
Gp3_im_re_a1 0 x3_im_a1 x3_re_a1 0 -262327540913.7152
Rp3_im_im_a1 0 x3_im_a1 6.71721917054064e-11
Cx4_re_a1 x4_re_a1 0 1.0
Gx4_re_a1 0 x4_re_a1 p1 0 0.1414213562373095
Fx4_re_a1 0 x4_re_a1 V1 7.0710678118654755
Rp4_re_re_a1 0 x4_re_a1 6.373089120988855e-11
Gp4_re_im_a1 0 x4_re_a1 x4_im_a1 0 218318096813.21487
Cx4_im_a1 x4_im_a1 0 1.0
Gp4_im_re_a1 0 x4_im_a1 x4_re_a1 0 -218318096813.21487
Rp4_im_im_a1 0 x4_im_a1 6.373089120988855e-11
Cx5_re_a1 x5_re_a1 0 1.0
Gx5_re_a1 0 x5_re_a1 p1 0 0.1414213562373095
Fx5_re_a1 0 x5_re_a1 V1 7.0710678118654755
Rp5_re_re_a1 0 x5_re_a1 6.440861041643573e-11
Gp5_re_im_a1 0 x5_re_a1 x5_im_a1 0 174592015736.0517
Cx5_im_a1 x5_im_a1 0 1.0
Gp5_im_re_a1 0 x5_im_a1 x5_re_a1 0 -174592015736.0517
Rp5_im_im_a1 0 x5_im_a1 6.440861041643573e-11
Cx6_re_a1 x6_re_a1 0 1.0
Gx6_re_a1 0 x6_re_a1 p1 0 0.1414213562373095
Fx6_re_a1 0 x6_re_a1 V1 7.0710678118654755
Rp6_re_re_a1 0 x6_re_a1 6.53938629165566e-11
Gp6_re_im_a1 0 x6_re_a1 x6_im_a1 0 130889967614.0941
Cx6_im_a1 x6_im_a1 0 1.0
Gp6_im_re_a1 0 x6_im_a1 x6_re_a1 0 -130889967614.0941
Rp6_im_im_a1 0 x6_im_a1 6.53938629165566e-11
Cx7_re_a1 x7_re_a1 0 1.0
Gx7_re_a1 0 x7_re_a1 p1 0 0.1414213562373095
Fx7_re_a1 0 x7_re_a1 V1 7.0710678118654755
Rp7_re_re_a1 0 x7_re_a1 6.659131890324554e-11
Gp7_re_im_a1 0 x7_re_a1 x7_im_a1 0 87152219067.44771
Cx7_im_a1 x7_im_a1 0 1.0
Gp7_im_re_a1 0 x7_im_a1 x7_re_a1 0 -87152219067.44771
Rp7_im_im_a1 0 x7_im_a1 6.659131890324554e-11
Cx8_re_a1 x8_re_a1 0 1.0
Gx8_re_a1 0 x8_re_a1 p1 0 0.1414213562373095
Fx8_re_a1 0 x8_re_a1 V1 7.0710678118654755
Rp8_re_re_a1 0 x8_re_a1 6.776175054208851e-11
Gp8_re_im_a1 0 x8_re_a1 x8_im_a1 0 43381529970.948
Cx8_im_a1 x8_im_a1 0 1.0
Gp8_im_re_a1 0 x8_im_a1 x8_re_a1 0 -43381529970.948
Rp8_im_im_a1 0 x8_im_a1 6.776175054208851e-11
Cx9_a1 x9_a1 0 1.0
Gx9_a1 0 x9_a1 p1 0 0.07071067811865475
Fx9_a1 0 x9_a1 V1 3.5355339059327378
Rp9_a1 0 x9_a1 6.778729912468209e-11
Cx10_re_a1 x10_re_a1 0 1.0
Gx10_re_a1 0 x10_re_a1 p1 0 0.1414213562373095
Fx10_re_a1 0 x10_re_a1 V1 7.0710678118654755
Rp10_re_re_a1 0 x10_re_a1 5.266227603617706e-10
Gp10_re_im_a1 0 x10_re_a1 x10_im_a1 0 2228171539.324897
Cx10_im_a1 x10_im_a1 0 1.0
Gp10_im_re_a1 0 x10_im_a1 x10_re_a1 0 -2228171539.324897
Rp10_im_im_a1 0 x10_im_a1 5.266227603617706e-10
Cx11_a1 x11_a1 0 1.0
Gx11_a1 0 x11_a1 p1 0 0.07071067811865475
Fx11_a1 0 x11_a1 V1 3.5355339059327378
Rp11_a1 0 x11_a1 5.172809035131532e-10
*
* Port network for port 2
V2 p2 s2 0
R2 s2 0 50.0
Gd2_1 0 s2 p1 0 -0.0016856930057705024
Fd2_1 0 s2 V1 -0.08428465028852512
Gr1_2_1 0 s2 x1_a1 0 114980691786.52333
Gr2_re_2_1 0 s2 x2_re_a1 0 -3439807808.414713
Gr2_im_2_1 0 s2 x2_im_a1 0 2514561760.7022943
Gr3_re_2_1 0 s2 x3_re_a1 0 4423321369.533221
Gr3_im_2_1 0 s2 x3_im_a1 0 -651374200.6221441
Gr4_re_2_1 0 s2 x4_re_a1 0 -4684893909.527277
Gr4_im_2_1 0 s2 x4_im_a1 0 -61217124.355229184
Gr5_re_2_1 0 s2 x5_re_a1 0 4712777508.873271
Gr5_im_2_1 0 s2 x5_im_a1 0 73744102.59193528
Gr6_re_2_1 0 s2 x6_re_a1 0 -4702204173.996919
Gr6_im_2_1 0 s2 x6_im_a1 0 -68486113.0385877
Gr7_re_2_1 0 s2 x7_re_a1 0 4691734541.675553
Gr7_im_2_1 0 s2 x7_im_a1 0 92677089.01510254
Gr8_re_2_1 0 s2 x8_re_a1 0 -4725312491.317949
Gr8_im_2_1 0 s2 x8_im_a1 0 -120007193.34835534
Gr9_2_1 0 s2 x9_a1 0 4665975028.099111
Gr10_re_2_1 0 s2 x10_re_a1 0 -560743.6183148772
Gr10_im_2_1 0 s2 x10_im_a1 0 2135652.8297383706
Gr11_2_1 0 s2 x11_a1 0 -1099763.155693093
Gd2_2 0 s2 p2 0 -0.05599437861010728
Fd2_2 0 s2 V2 -2.7997189305053642
Gr1_2_2 0 s2 x1_a2 0 3749671826091.7417
Gr2_re_2_2 0 s2 x2_re_a2 0 -20119730888.36094
Gr2_im_2_2 0 s2 x2_im_a2 0 -7615793267.563459
Gr3_re_2_2 0 s2 x3_re_a2 0 -4582270774.515796
Gr3_im_2_2 0 s2 x3_im_a2 0 327605610.7607822
Gr4_re_2_2 0 s2 x4_re_a2 0 -4687608450.879956
Gr4_im_2_2 0 s2 x4_im_a2 0 -60815242.74458649
Gr5_re_2_2 0 s2 x5_re_a2 0 -4703207822.656032
Gr5_im_2_2 0 s2 x5_im_a2 0 -73675770.72488862
Gr6_re_2_2 0 s2 x6_re_a2 0 -4696210203.282378
Gr6_im_2_2 0 s2 x6_im_a2 0 -70184505.1691104
Gr7_re_2_2 0 s2 x7_re_a2 0 -4690028374.353796
Gr7_im_2_2 0 s2 x7_im_a2 0 -82816399.82581523
Gr8_re_2_2 0 s2 x8_re_a2 0 -4721421341.403382
Gr8_im_2_2 0 s2 x8_im_a2 0 -106419878.93335322
Gr9_2_2 0 s2 x9_a2 0 -4689776981.430431
Gr10_re_2_2 0 s2 x10_re_a2 0 1043910.4473997038
Gr10_im_2_2 0 s2 x10_im_a2 0 -118841.77270125736
Gr11_2_2 0 s2 x11_a2 0 4592739.718917729
*
* State networks driven by port 2
Cx1_a2 x1_a2 0 1.0
Gx1_a2 0 x1_a2 p2 0 0.07071067811865475
Fx1_a2 0 x1_a2 V2 3.5355339059327378
Rp1_a2 0 x1_a2 3.1658774695127977e-13
Cx2_re_a2 x2_re_a2 0 1.0
Gx2_re_a2 0 x2_re_a2 p2 0 0.1414213562373095
Fx2_re_a2 0 x2_re_a2 V2 7.0710678118654755
Rp2_re_re_a2 0 x2_re_a2 3.094780737837525e-11
Gp2_re_im_a2 0 x2_re_a2 x2_im_a2 0 338816889165.91437
Cx2_im_a2 x2_im_a2 0 1.0
Gp2_im_re_a2 0 x2_im_a2 x2_re_a2 0 -338816889165.91437
Rp2_im_im_a2 0 x2_im_a2 3.094780737837525e-11
Cx3_re_a2 x3_re_a2 0 1.0
Gx3_re_a2 0 x3_re_a2 p2 0 0.1414213562373095
Fx3_re_a2 0 x3_re_a2 V2 7.0710678118654755
Rp3_re_re_a2 0 x3_re_a2 6.71721917054064e-11
Gp3_re_im_a2 0 x3_re_a2 x3_im_a2 0 262327540913.7152
Cx3_im_a2 x3_im_a2 0 1.0
Gp3_im_re_a2 0 x3_im_a2 x3_re_a2 0 -262327540913.7152
Rp3_im_im_a2 0 x3_im_a2 6.71721917054064e-11
Cx4_re_a2 x4_re_a2 0 1.0
Gx4_re_a2 0 x4_re_a2 p2 0 0.1414213562373095
Fx4_re_a2 0 x4_re_a2 V2 7.0710678118654755
Rp4_re_re_a2 0 x4_re_a2 6.373089120988855e-11
Gp4_re_im_a2 0 x4_re_a2 x4_im_a2 0 218318096813.21487
Cx4_im_a2 x4_im_a2 0 1.0
Gp4_im_re_a2 0 x4_im_a2 x4_re_a2 0 -218318096813.21487
Rp4_im_im_a2 0 x4_im_a2 6.373089120988855e-11
Cx5_re_a2 x5_re_a2 0 1.0
Gx5_re_a2 0 x5_re_a2 p2 0 0.1414213562373095
Fx5_re_a2 0 x5_re_a2 V2 7.0710678118654755
Rp5_re_re_a2 0 x5_re_a2 6.440861041643573e-11
Gp5_re_im_a2 0 x5_re_a2 x5_im_a2 0 174592015736.0517
Cx5_im_a2 x5_im_a2 0 1.0
Gp5_im_re_a2 0 x5_im_a2 x5_re_a2 0 -174592015736.0517
Rp5_im_im_a2 0 x5_im_a2 6.440861041643573e-11
Cx6_re_a2 x6_re_a2 0 1.0
Gx6_re_a2 0 x6_re_a2 p2 0 0.1414213562373095
Fx6_re_a2 0 x6_re_a2 V2 7.0710678118654755
Rp6_re_re_a2 0 x6_re_a2 6.53938629165566e-11
Gp6_re_im_a2 0 x6_re_a2 x6_im_a2 0 130889967614.0941
Cx6_im_a2 x6_im_a2 0 1.0
Gp6_im_re_a2 0 x6_im_a2 x6_re_a2 0 -130889967614.0941
Rp6_im_im_a2 0 x6_im_a2 6.53938629165566e-11
Cx7_re_a2 x7_re_a2 0 1.0
Gx7_re_a2 0 x7_re_a2 p2 0 0.1414213562373095
Fx7_re_a2 0 x7_re_a2 V2 7.0710678118654755
Rp7_re_re_a2 0 x7_re_a2 6.659131890324554e-11
Gp7_re_im_a2 0 x7_re_a2 x7_im_a2 0 87152219067.44771
Cx7_im_a2 x7_im_a2 0 1.0
Gp7_im_re_a2 0 x7_im_a2 x7_re_a2 0 -87152219067.44771
Rp7_im_im_a2 0 x7_im_a2 6.659131890324554e-11
Cx8_re_a2 x8_re_a2 0 1.0
Gx8_re_a2 0 x8_re_a2 p2 0 0.1414213562373095
Fx8_re_a2 0 x8_re_a2 V2 7.0710678118654755
Rp8_re_re_a2 0 x8_re_a2 6.776175054208851e-11
Gp8_re_im_a2 0 x8_re_a2 x8_im_a2 0 43381529970.948
Cx8_im_a2 x8_im_a2 0 1.0
Gp8_im_re_a2 0 x8_im_a2 x8_re_a2 0 -43381529970.948
Rp8_im_im_a2 0 x8_im_a2 6.776175054208851e-11
Cx9_a2 x9_a2 0 1.0
Gx9_a2 0 x9_a2 p2 0 0.07071067811865475
Fx9_a2 0 x9_a2 V2 3.5355339059327378
Rp9_a2 0 x9_a2 6.778729912468209e-11
Cx10_re_a2 x10_re_a2 0 1.0
Gx10_re_a2 0 x10_re_a2 p2 0 0.1414213562373095
Fx10_re_a2 0 x10_re_a2 V2 7.0710678118654755
Rp10_re_re_a2 0 x10_re_a2 5.266227603617706e-10
Gp10_re_im_a2 0 x10_re_a2 x10_im_a2 0 2228171539.324897
Cx10_im_a2 x10_im_a2 0 1.0
Gp10_im_re_a2 0 x10_im_a2 x10_re_a2 0 -2228171539.324897
Rp10_im_im_a2 0 x10_im_a2 5.266227603617706e-10
Cx11_a2 x11_a2 0 1.0
Gx11_a2 0 x11_a2 p2 0 0.07071067811865475
Fx11_a2 0 x11_a2 V2 3.5355339059327378
Rp11_a2 0 x11_a2 5.172809035131532e-10
.ENDS s_equivalent
