* EQUIVALENT CIRCUIT FOR VECTOR FITTED S-MATRIX
* Created using scikit-rf vectorFitting.py
*
.SUBCKT s_equivalent p1 p2 p3 p4
*
* Port network for port 1
V1 p1 s1 0
R1 s1 0 50.0
Gd1_1 0 s1 p1 0 7.260681220548722e-05
Fd1_1 0 s1 V1 0.003630340610274361
Gr1_re_1_1 0 s1 x1_re_a1 0 -33001167.305772625
Gr1_im_1_1 0 s1 x1_im_a1 0 -2957399390.3025904
Gr2_re_1_1 0 s1 x2_re_a1 0 23232754336.912304
Gr2_im_1_1 0 s1 x2_im_a1 0 -2202713522.214869
Gr3_re_1_1 0 s1 x3_re_a1 0 -34826972004.73593
Gr3_im_1_1 0 s1 x3_im_a1 0 -20708516859.57584
Gr4_1_1 0 s1 x4_a1 0 -4343296.185547169
Gr5_re_1_1 0 s1 x5_re_a1 0 -6527419318.687704
Gr5_im_1_1 0 s1 x5_im_a1 0 -717060043.7535005
Gr6_1_1 0 s1 x6_a1 0 3545218768.092161
Gd1_2 0 s1 p2 0 0.0057196677476184545
Fd1_2 0 s1 V2 0.28598338738092277
Gr1_re_1_2 0 s1 x1_re_a2 0 9247587503.580122
Gr1_im_1_2 0 s1 x1_im_a2 0 -14075193379.369188
Gr2_re_1_2 0 s1 x2_re_a2 0 -7449453507.136441
Gr2_im_1_2 0 s1 x2_im_a2 0 15547790295.17895
Gr3_re_1_2 0 s1 x3_re_a2 0 -9021213110.400026
Gr3_im_1_2 0 s1 x3_im_a2 0 -51236154436.92843
Gr4_1_2 0 s1 x4_a2 0 -163180.73853699793
Gr5_re_1_2 0 s1 x5_re_a2 0 -4798682368.092117
Gr5_im_1_2 0 s1 x5_im_a2 0 13736227502.67451
Gr6_1_2 0 s1 x6_a2 0 -19402763389.46812
Gd1_3 0 s1 p3 0 -0.00036438972112726035
Fd1_3 0 s1 V3 -0.01821948605636302
Gr1_re_1_3 0 s1 x1_re_a3 0 31916716269.93498
Gr1_im_1_3 0 s1 x1_im_a3 0 19112583812.25881
Gr2_re_1_3 0 s1 x2_re_a3 0 -13222217549.663137
Gr2_im_1_3 0 s1 x2_im_a3 0 17665377867.817253
Gr3_re_1_3 0 s1 x3_re_a3 0 -33951594462.02287
Gr3_im_1_3 0 s1 x3_im_a3 0 -43196866815.111916
Gr4_1_3 0 s1 x4_a3 0 4275274.667179357
Gr5_re_1_3 0 s1 x5_re_a3 0 12353559393.182465
Gr5_im_1_3 0 s1 x5_im_a3 0 -11435841939.212122
Gr6_1_3 0 s1 x6_a3 0 23917418107.687046
Gd1_4 0 s1 p4 0 5.780283412748834e-05
Fd1_4 0 s1 V4 0.002890141706374417
Gr1_re_1_4 0 s1 x1_re_a4 0 19283581881.002167
Gr1_im_1_4 0 s1 x1_im_a4 0 -8177164502.926022
Gr2_re_1_4 0 s1 x2_re_a4 0 20580394858.47782
Gr2_im_1_4 0 s1 x2_im_a4 0 -3518176965.227322
Gr3_re_1_4 0 s1 x3_re_a4 0 -46278688249.63373
Gr3_im_1_4 0 s1 x3_im_a4 0 -19844211067.644432
Gr4_1_4 0 s1 x4_a4 0 5030763.950512429
Gr5_re_1_4 0 s1 x5_re_a4 0 1154585999.101908
Gr5_im_1_4 0 s1 x5_im_a4 0 -4853296965.161308
Gr6_1_4 0 s1 x6_a4 0 -8425501453.112738
*
* State networks driven by port 1
Cx1_re_a1 x1_re_a1 0 1.0
Gx1_re_a1 0 x1_re_a1 p1 0 0.1414213562373095
Fx1_re_a1 0 x1_re_a1 V1 7.0710678118654755
Rp1_re_re_a1 0 x1_re_a1 7.265956860616756e-12
Gp1_re_im_a1 0 x1_re_a1 x1_im_a1 0 572815983367.4526
Cx1_im_a1 x1_im_a1 0 1.0
Gp1_im_re_a1 0 x1_im_a1 x1_re_a1 0 -572815983367.4526
Rp1_im_im_a1 0 x1_im_a1 7.265956860616756e-12
Cx2_re_a1 x2_re_a1 0 1.0
Gx2_re_a1 0 x2_re_a1 p1 0 0.1414213562373095
Fx2_re_a1 0 x2_re_a1 V1 7.0710678118654755
Rp2_re_re_a1 0 x2_re_a1 6.803467392229221e-12
Gp2_re_im_a1 0 x2_re_a1 x2_im_a1 0 395441498330.00323
Cx2_im_a1 x2_im_a1 0 1.0
Gp2_im_re_a1 0 x2_im_a1 x2_re_a1 0 -395441498330.00323
Rp2_im_im_a1 0 x2_im_a1 6.803467392229221e-12
Cx3_re_a1 x3_re_a1 0 1.0
Gx3_re_a1 0 x3_re_a1 p1 0 0.1414213562373095
Fx3_re_a1 0 x3_re_a1 V1 7.0710678118654755
Rp3_re_re_a1 0 x3_re_a1 4.614973865662602e-12
Gp3_re_im_a1 0 x3_re_a1 x3_im_a1 0 290216169888.9015
Cx3_im_a1 x3_im_a1 0 1.0
Gp3_im_re_a1 0 x3_im_a1 x3_re_a1 0 -290216169888.9015
Rp3_im_im_a1 0 x3_im_a1 4.614973865662602e-12
Cx4_a1 x4_a1 0 1.0
Gx4_a1 0 x4_a1 p1 0 0.07071067811865475
Fx4_a1 0 x4_a1 V1 3.5355339059327378
Rp4_a1 0 x4_a1 4.409490349112835e-11
Cx5_re_a1 x5_re_a1 0 1.0
Gx5_re_a1 0 x5_re_a1 p1 0 0.1414213562373095
Fx5_re_a1 0 x5_re_a1 V1 7.0710678118654755
Rp5_re_re_a1 0 x5_re_a1 5.944748916473448e-12
Gp5_re_im_a1 0 x5_re_a1 x5_im_a1 0 77979147588.22144
Cx5_im_a1 x5_im_a1 0 1.0
Gp5_im_re_a1 0 x5_im_a1 x5_re_a1 0 -77979147588.22144
Rp5_im_im_a1 0 x5_im_a1 5.944748916473448e-12
Cx6_a1 x6_a1 0 1.0
Gx6_a1 0 x6_a1 p1 0 0.07071067811865475
Fx6_a1 0 x6_a1 V1 3.5355339059327378
Rp6_a1 0 x6_a1 7.259790773231773e-12
*
* Port network for port 2
V2 p2 s2 0
R2 s2 0 50.0
Gd2_1 0 s2 p1 0 0.005719667747678166
Fd2_1 0 s2 V1 0.2859833873839083
Gr1_re_2_1 0 s2 x1_re_a1 0 9247587503.533278
Gr1_im_2_1 0 s2 x1_im_a1 0 -14075193379.63031
Gr2_re_2_1 0 s2 x2_re_a1 0 -7449453507.225638
Gr2_im_2_1 0 s2 x2_im_a1 0 15547790295.359089
Gr3_re_2_1 0 s2 x3_re_a1 0 -9021213110.50428
Gr3_im_2_1 0 s2 x3_im_a1 0 -51236154437.28675
Gr4_2_1 0 s2 x4_a1 0 -163180.7378577855
Gr5_re_2_1 0 s2 x5_re_a1 0 -4798682368.182566
Gr5_im_2_1 0 s2 x5_im_a1 0 13736227502.637674
Gr6_2_1 0 s2 x6_a1 0 -19402763389.64742
Gd2_2 0 s2 p2 0 7.260681221175617e-05
Fd2_2 0 s2 V2 0.003630340610587809
Gr1_re_2_2 0 s2 x1_re_a2 0 -33001167.309350353
Gr1_im_2_2 0 s2 x1_im_a2 0 -2957399390.3302755
Gr2_re_2_2 0 s2 x2_re_a2 0 23232754336.902035
Gr2_im_2_2 0 s2 x2_im_a2 0 -2202713522.1873837
Gr3_re_2_2 0 s2 x3_re_a2 0 -34826972004.7422
Gr3_im_2_2 0 s2 x3_im_a2 0 -20708516859.624924
Gr4_2_2 0 s2 x4_a2 0 -4343296.185485327
Gr5_re_2_2 0 s2 x5_re_a2 0 -6527419318.695952
Gr5_im_2_2 0 s2 x5_im_a2 0 -717060043.7536246
Gr6_2_2 0 s2 x6_a2 0 3545218768.070206
Gd2_3 0 s2 p3 0 5.7802834111114535e-05
Fd2_3 0 s2 V3 0.002890141705555727
Gr1_re_2_3 0 s2 x1_re_a3 0 19283581880.877766
Gr1_im_2_3 0 s2 x1_im_a3 0 -8177164502.541969
Gr2_re_2_3 0 s2 x2_re_a3 0 20580394858.500988
Gr2_im_2_3 0 s2 x2_im_a3 0 -3518176965.3465223
Gr3_re_2_3 0 s2 x3_re_a3 0 -46278688249.35856
Gr3_im_2_3 0 s2 x3_im_a3 0 -19844211067.713722
Gr4_2_3 0 s2 x4_a3 0 5030763.949918692
Gr5_re_2_3 0 s2 x5_re_a3 0 1154585999.1582081
Gr5_im_2_3 0 s2 x5_im_a3 0 -4853296965.056045
Gr6_2_3 0 s2 x6_a3 0 -8425501453.141163
Gd2_4 0 s2 p4 0 -0.00036438972112836537
Fd2_4 0 s2 V4 -0.01821948605641827
Gr1_re_2_4 0 s2 x1_re_a4 0 31916716269.919212
Gr1_im_2_4 0 s2 x1_im_a4 0 19112583812.302013
Gr2_re_2_4 0 s2 x2_re_a4 0 -13222217549.659496
Gr2_im_2_4 0 s2 x2_im_a4 0 17665377867.79988
Gr3_re_2_4 0 s2 x3_re_a4 0 -33951594461.99641
Gr3_im_2_4 0 s2 x3_im_a4 0 -43196866815.120384
Gr4_2_4 0 s2 x4_a4 0 4275274.667107617
Gr5_re_2_4 0 s2 x5_re_a4 0 12353559393.188238
Gr5_im_2_4 0 s2 x5_im_a4 0 -11435841939.19952
Gr6_2_4 0 s2 x6_a4 0 23917418107.68269
*
* State networks driven by port 2
Cx1_re_a2 x1_re_a2 0 1.0
Gx1_re_a2 0 x1_re_a2 p2 0 0.1414213562373095
Fx1_re_a2 0 x1_re_a2 V2 7.0710678118654755
Rp1_re_re_a2 0 x1_re_a2 7.265956860616756e-12
Gp1_re_im_a2 0 x1_re_a2 x1_im_a2 0 572815983367.4526
Cx1_im_a2 x1_im_a2 0 1.0
Gp1_im_re_a2 0 x1_im_a2 x1_re_a2 0 -572815983367.4526
Rp1_im_im_a2 0 x1_im_a2 7.265956860616756e-12
Cx2_re_a2 x2_re_a2 0 1.0
Gx2_re_a2 0 x2_re_a2 p2 0 0.1414213562373095
Fx2_re_a2 0 x2_re_a2 V2 7.0710678118654755
Rp2_re_re_a2 0 x2_re_a2 6.803467392229221e-12
Gp2_re_im_a2 0 x2_re_a2 x2_im_a2 0 395441498330.00323
Cx2_im_a2 x2_im_a2 0 1.0
Gp2_im_re_a2 0 x2_im_a2 x2_re_a2 0 -395441498330.00323
Rp2_im_im_a2 0 x2_im_a2 6.803467392229221e-12
Cx3_re_a2 x3_re_a2 0 1.0
Gx3_re_a2 0 x3_re_a2 p2 0 0.1414213562373095
Fx3_re_a2 0 x3_re_a2 V2 7.0710678118654755
Rp3_re_re_a2 0 x3_re_a2 4.614973865662602e-12
Gp3_re_im_a2 0 x3_re_a2 x3_im_a2 0 290216169888.9015
Cx3_im_a2 x3_im_a2 0 1.0
Gp3_im_re_a2 0 x3_im_a2 x3_re_a2 0 -290216169888.9015
Rp3_im_im_a2 0 x3_im_a2 4.614973865662602e-12
Cx4_a2 x4_a2 0 1.0
Gx4_a2 0 x4_a2 p2 0 0.07071067811865475
Fx4_a2 0 x4_a2 V2 3.5355339059327378
Rp4_a2 0 x4_a2 4.409490349112835e-11
Cx5_re_a2 x5_re_a2 0 1.0
Gx5_re_a2 0 x5_re_a2 p2 0 0.1414213562373095
Fx5_re_a2 0 x5_re_a2 V2 7.0710678118654755
Rp5_re_re_a2 0 x5_re_a2 5.944748916473448e-12
Gp5_re_im_a2 0 x5_re_a2 x5_im_a2 0 77979147588.22144
Cx5_im_a2 x5_im_a2 0 1.0
Gp5_im_re_a2 0 x5_im_a2 x5_re_a2 0 -77979147588.22144
Rp5_im_im_a2 0 x5_im_a2 5.944748916473448e-12
Cx6_a2 x6_a2 0 1.0
Gx6_a2 0 x6_a2 p2 0 0.07071067811865475
Fx6_a2 0 x6_a2 V2 3.5355339059327378
Rp6_a2 0 x6_a2 7.259790773231773e-12
*
* Port network for port 3
V3 p3 s3 0
R3 s3 0 50.0
Gd3_1 0 s3 p1 0 -0.0003643897211272926
Fd3_1 0 s3 V1 -0.01821948605636463
Gr1_re_3_1 0 s3 x1_re_a1 0 31916716269.934982
Gr1_im_3_1 0 s3 x1_im_a1 0 19112583812.258743
Gr2_re_3_1 0 s3 x2_re_a1 0 -13222217549.663368
Gr2_im_3_1 0 s3 x2_im_a1 0 17665377867.8173
Gr3_re_3_1 0 s3 x3_re_a1 0 -33951594462.02271
Gr3_im_3_1 0 s3 x3_im_a1 0 -43196866815.11153
Gr4_3_1 0 s3 x4_a1 0 4275274.6671807105
Gr5_re_3_1 0 s3 x5_re_a1 0 12353559393.18257
Gr5_im_3_1 0 s3 x5_im_a1 0 -11435841939.211702
Gr6_3_1 0 s3 x6_a1 0 23917418107.687443
Gd3_2 0 s3 p2 0 5.7802834127548865e-05
Fd3_2 0 s3 V2 0.0028901417063774437
Gr1_re_3_2 0 s3 x1_re_a2 0 19283581881.002155
Gr1_im_3_2 0 s3 x1_im_a2 0 -8177164502.926152
Gr2_re_3_2 0 s3 x2_re_a2 0 20580394858.47792
Gr2_im_3_2 0 s3 x2_im_a2 0 -3518176965.227379
Gr3_re_3_2 0 s3 x3_re_a2 0 -46278688249.63399
Gr3_im_3_2 0 s3 x3_im_a2 0 -19844211067.644844
Gr4_3_2 0 s3 x4_a2 0 5030763.950513486
Gr5_re_3_2 0 s3 x5_re_a2 0 1154585999.1017227
Gr5_im_3_2 0 s3 x5_im_a2 0 -4853296965.161742
Gr6_3_2 0 s3 x6_a2 0 -8425501453.113133
Gd3_3 0 s3 p3 0 7.260681220538501e-05
Fd3_3 0 s3 V3 0.0036303406102692506
Gr1_re_3_3 0 s3 x1_re_a3 0 -33001167.305888858
Gr1_im_3_3 0 s3 x1_im_a3 0 -2957399390.3020854
Gr2_re_3_3 0 s3 x2_re_a3 0 23232754336.912346
Gr2_im_3_3 0 s3 x2_im_a3 0 -2202713522.2145123
Gr3_re_3_3 0 s3 x3_re_a3 0 -34826972004.73513
Gr3_im_3_3 0 s3 x3_im_a3 0 -20708516859.575645
Gr4_3_3 0 s3 x4_a3 0 -4343296.185547471
Gr5_re_3_3 0 s3 x5_re_a3 0 -6527419318.68742
Gr5_im_3_3 0 s3 x5_im_a3 0 -717060043.7533048
Gr6_3_3 0 s3 x6_a3 0 3545218768.092295
Gd3_4 0 s3 p4 0 0.005719667747618475
Fd3_4 0 s3 V4 0.28598338738092377
Gr1_re_3_4 0 s3 x1_re_a4 0 9247587503.580042
Gr1_im_3_4 0 s3 x1_im_a4 0 -14075193379.369085
Gr2_re_3_4 0 s3 x2_re_a4 0 -7449453507.136288
Gr2_im_3_4 0 s3 x2_im_a4 0 15547790295.179037
Gr3_re_3_4 0 s3 x3_re_a4 0 -9021213110.400013
Gr3_im_3_4 0 s3 x3_im_a4 0 -51236154436.92877
Gr4_3_4 0 s3 x4_a4 0 -163180.73853656292
Gr5_re_3_4 0 s3 x5_re_a4 0 -4798682368.092214
Gr5_im_3_4 0 s3 x5_im_a4 0 13736227502.674288
Gr6_3_4 0 s3 x6_a4 0 -19402763389.46832
*
* State networks driven by port 3
Cx1_re_a3 x1_re_a3 0 1.0
Gx1_re_a3 0 x1_re_a3 p3 0 0.1414213562373095
Fx1_re_a3 0 x1_re_a3 V3 7.0710678118654755
Rp1_re_re_a3 0 x1_re_a3 7.265956860616756e-12
Gp1_re_im_a3 0 x1_re_a3 x1_im_a3 0 572815983367.4526
Cx1_im_a3 x1_im_a3 0 1.0
Gp1_im_re_a3 0 x1_im_a3 x1_re_a3 0 -572815983367.4526
Rp1_im_im_a3 0 x1_im_a3 7.265956860616756e-12
Cx2_re_a3 x2_re_a3 0 1.0
Gx2_re_a3 0 x2_re_a3 p3 0 0.1414213562373095
Fx2_re_a3 0 x2_re_a3 V3 7.0710678118654755
Rp2_re_re_a3 0 x2_re_a3 6.803467392229221e-12
Gp2_re_im_a3 0 x2_re_a3 x2_im_a3 0 395441498330.00323
Cx2_im_a3 x2_im_a3 0 1.0
Gp2_im_re_a3 0 x2_im_a3 x2_re_a3 0 -395441498330.00323
Rp2_im_im_a3 0 x2_im_a3 6.803467392229221e-12
Cx3_re_a3 x3_re_a3 0 1.0
Gx3_re_a3 0 x3_re_a3 p3 0 0.1414213562373095
Fx3_re_a3 0 x3_re_a3 V3 7.0710678118654755
Rp3_re_re_a3 0 x3_re_a3 4.614973865662602e-12
Gp3_re_im_a3 0 x3_re_a3 x3_im_a3 0 290216169888.9015
Cx3_im_a3 x3_im_a3 0 1.0
Gp3_im_re_a3 0 x3_im_a3 x3_re_a3 0 -290216169888.9015
Rp3_im_im_a3 0 x3_im_a3 4.614973865662602e-12
Cx4_a3 x4_a3 0 1.0
Gx4_a3 0 x4_a3 p3 0 0.07071067811865475
Fx4_a3 0 x4_a3 V3 3.5355339059327378
Rp4_a3 0 x4_a3 4.409490349112835e-11
Cx5_re_a3 x5_re_a3 0 1.0
Gx5_re_a3 0 x5_re_a3 p3 0 0.1414213562373095
Fx5_re_a3 0 x5_re_a3 V3 7.0710678118654755
Rp5_re_re_a3 0 x5_re_a3 5.944748916473448e-12
Gp5_re_im_a3 0 x5_re_a3 x5_im_a3 0 77979147588.22144
Cx5_im_a3 x5_im_a3 0 1.0
Gp5_im_re_a3 0 x5_im_a3 x5_re_a3 0 -77979147588.22144
Rp5_im_im_a3 0 x5_im_a3 5.944748916473448e-12
Cx6_a3 x6_a3 0 1.0
Gx6_a3 0 x6_a3 p3 0 0.07071067811865475
Fx6_a3 0 x6_a3 V3 3.5355339059327378
Rp6_a3 0 x6_a3 7.259790773231773e-12
*
* Port network for port 4
V4 p4 s4 0
R4 s4 0 50.0
Gd4_1 0 s4 p1 0 5.780283411111286e-05
Fd4_1 0 s4 V1 0.002890141705555643
Gr1_re_4_1 0 s4 x1_re_a1 0 19283581880.87762
Gr1_im_4_1 0 s4 x1_im_a1 0 -8177164502.542051
Gr2_re_4_1 0 s4 x2_re_a1 0 20580394858.50078
Gr2_im_4_1 0 s4 x2_im_a1 0 -3518176965.3464637
Gr3_re_4_1 0 s4 x3_re_a1 0 -46278688249.35841
Gr3_im_4_1 0 s4 x3_im_a1 0 -19844211067.713257
Gr4_4_1 0 s4 x4_a1 0 5030763.949914365
Gr5_re_4_1 0 s4 x5_re_a1 0 1154585999.158316
Gr5_im_4_1 0 s4 x5_im_a1 0 -4853296965.055621
Gr6_4_1 0 s4 x6_a1 0 -8425501453.140755
Gd4_2 0 s4 p2 0 -0.00036438972112832075
Fd4_2 0 s4 V2 -0.01821948605641604
Gr1_re_4_2 0 s4 x1_re_a2 0 31916716269.919468
Gr1_im_4_2 0 s4 x1_im_a2 0 19112583812.302048
Gr2_re_4_2 0 s4 x2_re_a2 0 -13222217549.659124
Gr2_im_4_2 0 s4 x2_im_a2 0 17665377867.799717
Gr3_re_4_2 0 s4 x3_re_a2 0 -33951594461.99677
Gr3_im_4_2 0 s4 x3_im_a2 0 -43196866815.12139
Gr4_4_2 0 s4 x4_a2 0 4275274.667112257
Gr5_re_4_2 0 s4 x5_re_a2 0 12353559393.187944
Gr5_im_4_2 0 s4 x5_im_a2 0 -11435841939.200636
Gr6_4_2 0 s4 x6_a2 0 23917418107.68162
Gd4_3 0 s4 p3 0 0.005719667747678187
Fd4_3 0 s4 V3 0.2859833873839094
Gr1_re_4_3 0 s4 x1_re_a3 0 9247587503.533293
Gr1_im_4_3 0 s4 x1_im_a3 0 -14075193379.630346
Gr2_re_4_3 0 s4 x2_re_a3 0 -7449453507.225509
Gr2_im_4_3 0 s4 x2_im_a3 0 15547790295.359081
Gr3_re_4_3 0 s4 x3_re_a3 0 -9021213110.50439
Gr3_im_4_3 0 s4 x3_im_a3 0 -51236154437.287094
Gr4_4_3 0 s4 x4_a3 0 -163180.7378562869
Gr5_re_4_3 0 s4 x5_re_a3 0 -4798682368.182669
Gr5_im_4_3 0 s4 x5_im_a3 0 13736227502.637306
Gr6_4_3 0 s4 x6_a3 0 -19402763389.647766
Gd4_4 0 s4 p4 0 7.260681221166249e-05
Fd4_4 0 s4 V4 0.003630340610583124
Gr1_re_4_4 0 s4 x1_re_a4 0 -33001167.309560817
Gr1_im_4_4 0 s4 x1_im_a4 0 -2957399390.329663
Gr2_re_4_4 0 s4 x2_re_a4 0 23232754336.902153
Gr2_im_4_4 0 s4 x2_im_a4 0 -2202713522.1870217
Gr3_re_4_4 0 s4 x3_re_a4 0 -34826972004.74154
Gr3_im_4_4 0 s4 x3_im_a4 0 -20708516859.62464
Gr4_4_4 0 s4 x4_a4 0 -4343296.185489472
Gr5_re_4_4 0 s4 x5_re_a4 0 -6527419318.69574
Gr5_im_4_4 0 s4 x5_im_a4 0 -717060043.7528973
Gr6_4_4 0 s4 x6_a4 0 3545218768.0709295
*
* State networks driven by port 4
Cx1_re_a4 x1_re_a4 0 1.0
Gx1_re_a4 0 x1_re_a4 p4 0 0.1414213562373095
Fx1_re_a4 0 x1_re_a4 V4 7.0710678118654755
Rp1_re_re_a4 0 x1_re_a4 7.265956860616756e-12
Gp1_re_im_a4 0 x1_re_a4 x1_im_a4 0 572815983367.4526
Cx1_im_a4 x1_im_a4 0 1.0
Gp1_im_re_a4 0 x1_im_a4 x1_re_a4 0 -572815983367.4526
Rp1_im_im_a4 0 x1_im_a4 7.265956860616756e-12
Cx2_re_a4 x2_re_a4 0 1.0
Gx2_re_a4 0 x2_re_a4 p4 0 0.1414213562373095
Fx2_re_a4 0 x2_re_a4 V4 7.0710678118654755
Rp2_re_re_a4 0 x2_re_a4 6.803467392229221e-12
Gp2_re_im_a4 0 x2_re_a4 x2_im_a4 0 395441498330.00323
Cx2_im_a4 x2_im_a4 0 1.0
Gp2_im_re_a4 0 x2_im_a4 x2_re_a4 0 -395441498330.00323
Rp2_im_im_a4 0 x2_im_a4 6.803467392229221e-12
Cx3_re_a4 x3_re_a4 0 1.0
Gx3_re_a4 0 x3_re_a4 p4 0 0.1414213562373095
Fx3_re_a4 0 x3_re_a4 V4 7.0710678118654755
Rp3_re_re_a4 0 x3_re_a4 4.614973865662602e-12
Gp3_re_im_a4 0 x3_re_a4 x3_im_a4 0 290216169888.9015
Cx3_im_a4 x3_im_a4 0 1.0
Gp3_im_re_a4 0 x3_im_a4 x3_re_a4 0 -290216169888.9015
Rp3_im_im_a4 0 x3_im_a4 4.614973865662602e-12
Cx4_a4 x4_a4 0 1.0
Gx4_a4 0 x4_a4 p4 0 0.07071067811865475
Fx4_a4 0 x4_a4 V4 3.5355339059327378
Rp4_a4 0 x4_a4 4.409490349112835e-11
Cx5_re_a4 x5_re_a4 0 1.0
Gx5_re_a4 0 x5_re_a4 p4 0 0.1414213562373095
Fx5_re_a4 0 x5_re_a4 V4 7.0710678118654755
Rp5_re_re_a4 0 x5_re_a4 5.944748916473448e-12
Gp5_re_im_a4 0 x5_re_a4 x5_im_a4 0 77979147588.22144
Cx5_im_a4 x5_im_a4 0 1.0
Gp5_im_re_a4 0 x5_im_a4 x5_re_a4 0 -77979147588.22144
Rp5_im_im_a4 0 x5_im_a4 5.944748916473448e-12
Cx6_a4 x6_a4 0 1.0
Gx6_a4 0 x6_a4 p4 0 0.07071067811865475
Fx6_a4 0 x6_a4 V4 3.5355339059327378
Rp6_a4 0 x6_a4 7.259790773231773e-12
.ENDS s_equivalent
