* EQUIVALENT CIRCUIT FOR VECTOR FITTED S-MATRIX
* Created using scikit-rf vectorFitting.py
*
.SUBCKT s_equivalent p1 p2 p3 p4
*
* Port network for port 1
V1 p1 s1 0
R1 s1 0 50.0
Gd1_1 0 s1 p1 0 -0.00018108907880570393
Fd1_1 0 s1 V1 -0.009054453940285197
Gr1_1_1 0 s1 x1_a1 0 21063934701.69753
Gr2_re_1_1 0 s1 x2_re_a1 0 -57060731756.96564
Gr2_im_1_1 0 s1 x2_im_a1 0 7979168490.9102125
Gr3_1_1 0 s1 x3_a1 0 -94899.57859888353
Gd1_2 0 s1 p2 0 0.00810284374224544
Fd1_2 0 s1 V2 0.405142187112272
Gr1_1_2 0 s1 x1_a2 0 -298221946013.7913
Gr2_re_1_2 0 s1 x2_re_a2 0 62098451306.1167
Gr2_im_1_2 0 s1 x2_im_a2 0 -56888227602.3583
Gr3_1_2 0 s1 x3_a2 0 -3856.82840762657
Gd1_3 0 s1 p3 0 0.00631619797022266
Fd1_3 0 s1 V3 0.31580989851113306
Gr1_1_3 0 s1 x1_a3 0 421506516899.1006
Gr2_re_1_3 0 s1 x2_re_a3 0 -203537941026.73022
Gr2_im_1_3 0 s1 x2_im_a3 0 26750767008.912296
Gr3_1_3 0 s1 x3_a3 0 122775.14604967424
Gd1_4 0 s1 p4 0 -0.0024298989639173017
Fd1_4 0 s1 V4 -0.12149494819586508
Gr1_1_4 0 s1 x1_a4 0 77669564285.70964
Gr2_re_1_4 0 s1 x2_re_a4 0 8430688711.169214
Gr2_im_1_4 0 s1 x2_im_a4 0 10166262929.424774
Gr3_1_4 0 s1 x3_a4 0 8197.399932350101
*
* State networks driven by port 1
Cx1_a1 x1_a1 0 1.0
Gx1_a1 0 x1_a1 p1 0 0.07071067811865475
Fx1_a1 0 x1_a1 V1 3.5355339059327378
Rp1_a1 0 x1_a1 5.282047205639696e-13
Cx2_re_a1 x2_re_a1 0 1.0
Gx2_re_a1 0 x2_re_a1 p1 0 0.1414213562373095
Fx2_re_a1 0 x2_re_a1 V1 7.0710678118654755
Rp2_re_re_a1 0 x2_re_a1 4.751370536275971e-12
Gp2_re_im_a1 0 x2_re_a1 x2_im_a1 0 2848279117741.6416
Cx2_im_a1 x2_im_a1 0 1.0
Gp2_im_re_a1 0 x2_im_a1 x2_re_a1 0 -2848279117741.6416
Rp2_im_im_a1 0 x2_im_a1 4.751370536275971e-12
Cx3_a1 x3_a1 0 1.0
Gx3_a1 0 x3_a1 p1 0 0.07071067811865475
Fx3_a1 0 x3_a1 V1 3.5355339059327378
Rp3_a1 0 x3_a1 3.5276330254138835e-10
*
* Port network for port 2
V2 p2 s2 0
R2 s2 0 50.0
Gd2_1 0 s2 p1 0 0.008084528805124893
Fd2_1 0 s2 V1 0.40422644025624466
Gr1_2_1 0 s2 x1_a1 0 -297448230648.91925
Gr2_re_2_1 0 s2 x2_re_a1 0 61822647521.427505
Gr2_im_2_1 0 s2 x2_im_a1 0 -56694287796.04822
Gr3_2_1 0 s2 x3_a1 0 -3849.268943595454
Gd2_2 0 s2 p2 0 0.003439029174894943
Fd2_2 0 s2 V2 0.17195145874474715
Gr1_2_2 0 s2 x1_a2 0 -130202809261.668
Gr2_re_2_2 0 s2 x2_re_a2 0 -7392709156.66481
Gr2_im_2_2 0 s2 x2_im_a2 0 -29462789592.235367
Gr3_2_2 0 s2 x3_a2 0 -113591.27365186867
Gd2_3 0 s2 p3 0 -0.002442414399063577
Fd2_3 0 s2 V3 -0.12212071995317884
Gr1_2_3 0 s2 x1_a3 0 78393861108.53021
Gr2_re_2_3 0 s2 x2_re_a3 0 8085377710.343883
Gr2_im_2_3 0 s2 x2_im_a3 0 10435145056.918648
Gr3_2_3 0 s2 x3_a3 0 8225.549809826112
Gd2_4 0 s2 p4 0 0.008189447288981511
Fd2_4 0 s2 V4 0.4094723644490756
Gr1_2_4 0 s2 x1_a4 0 306382530383.2505
Gr2_re_2_4 0 s2 x2_re_a4 0 -146369237910.8627
Gr2_im_2_4 0 s2 x2_im_a4 0 -18178093575.29191
Gr3_2_4 0 s2 x3_a4 0 99913.10743446814
*
* State networks driven by port 2
Cx1_a2 x1_a2 0 1.0
Gx1_a2 0 x1_a2 p2 0 0.07071067811865475
Fx1_a2 0 x1_a2 V2 3.5355339059327378
Rp1_a2 0 x1_a2 5.282047205639696e-13
Cx2_re_a2 x2_re_a2 0 1.0
Gx2_re_a2 0 x2_re_a2 p2 0 0.1414213562373095
Fx2_re_a2 0 x2_re_a2 V2 7.0710678118654755
Rp2_re_re_a2 0 x2_re_a2 4.751370536275971e-12
Gp2_re_im_a2 0 x2_re_a2 x2_im_a2 0 2848279117741.6416
Cx2_im_a2 x2_im_a2 0 1.0
Gp2_im_re_a2 0 x2_im_a2 x2_re_a2 0 -2848279117741.6416
Rp2_im_im_a2 0 x2_im_a2 4.751370536275971e-12
Cx3_a2 x3_a2 0 1.0
Gx3_a2 0 x3_a2 p2 0 0.07071067811865475
Fx3_a2 0 x3_a2 V2 3.5355339059327378
Rp3_a2 0 x3_a2 3.5276330254138835e-10
*
* Port network for port 3
V3 p3 s3 0
R3 s3 0 50.0
Gd3_1 0 s3 p1 0 0.006316197970229146
Fd3_1 0 s3 V1 0.3158098985114573
Gr1_3_1 0 s3 x1_a1 0 421506516899.0301
Gr2_re_3_1 0 s3 x2_re_a1 0 -203537941026.81732
Gr2_im_3_1 0 s3 x2_im_a1 0 26750767008.98413
Gr3_3_1 0 s3 x3_a1 0 122775.14608154458
Gd3_2 0 s3 p2 0 -0.0024298989639261735
Fd3_2 0 s3 V2 -0.12149494819630868
Gr1_3_2 0 s3 x1_a2 0 77669564285.79785
Gr2_re_3_2 0 s3 x2_re_a2 0 8430688711.28085
Gr2_im_3_2 0 s3 x2_im_a2 0 10166262929.319841
Gr3_3_2 0 s3 x3_a2 0 8197.39991114377
Gd3_3 0 s3 p3 0 -0.00018108907881045531
Fd3_3 0 s3 V3 -0.009054453940522766
Gr1_3_3 0 s3 x1_a3 0 21063934701.75017
Gr2_re_3_3 0 s3 x2_re_a3 0 -57060731756.901535
Gr2_im_3_3 0 s3 x2_im_a3 0 7979168490.858256
Gr3_3_3 0 s3 x3_a3 0 -94899.57862539361
Gd3_4 0 s3 p4 0 0.00810284374225894
Fd3_4 0 s3 V4 0.405142187112947
Gr1_3_4 0 s3 x1_a4 0 -298221946013.9257
Gr2_re_3_4 0 s3 x2_re_a4 0 62098451305.9472
Gr2_im_3_4 0 s3 x2_im_a4 0 -56888227602.198875
Gr3_3_4 0 s3 x3_a4 0 -3856.828376408068
*
* State networks driven by port 3
Cx1_a3 x1_a3 0 1.0
Gx1_a3 0 x1_a3 p3 0 0.07071067811865475
Fx1_a3 0 x1_a3 V3 3.5355339059327378
Rp1_a3 0 x1_a3 5.282047205639696e-13
Cx2_re_a3 x2_re_a3 0 1.0
Gx2_re_a3 0 x2_re_a3 p3 0 0.1414213562373095
Fx2_re_a3 0 x2_re_a3 V3 7.0710678118654755
Rp2_re_re_a3 0 x2_re_a3 4.751370536275971e-12
Gp2_re_im_a3 0 x2_re_a3 x2_im_a3 0 2848279117741.6416
Cx2_im_a3 x2_im_a3 0 1.0
Gp2_im_re_a3 0 x2_im_a3 x2_re_a3 0 -2848279117741.6416
Rp2_im_im_a3 0 x2_im_a3 4.751370536275971e-12
Cx3_a3 x3_a3 0 1.0
Gx3_a3 0 x3_a3 p3 0 0.07071067811865475
Fx3_a3 0 x3_a3 V3 3.5355339059327378
Rp3_a3 0 x3_a3 3.5276330254138835e-10
*
* Port network for port 4
V4 p4 s4 0
R4 s4 0 50.0
Gd4_1 0 s4 p1 0 -0.0024424143990475554
Fd4_1 0 s4 V1 -0.12212071995237778
Gr1_4_1 0 s4 x1_a1 0 78393861108.36604
Gr2_re_4_1 0 s4 x2_re_a1 0 8085377710.138838
Gr2_im_4_1 0 s4 x2_im_a1 0 10435145057.104315
Gr3_4_1 0 s4 x3_a1 0 8225.54985754036
Gd4_2 0 s4 p2 0 0.008189447288952106
Fd4_2 0 s4 V2 0.4094723644476054
Gr1_4_2 0 s4 x1_a2 0 306382530383.54346
Gr2_re_4_2 0 s4 x2_re_a2 0 -146369237910.49185
Gr2_im_4_2 0 s4 x2_im_a2 0 -18178093575.63932
Gr3_4_2 0 s4 x3_a2 0 99913.10737088392
Gd4_3 0 s4 p3 0 0.008084528805110595
Fd4_3 0 s4 V3 0.4042264402555298
Gr1_4_3 0 s4 x1_a3 0 -297448230648.77295
Gr2_re_4_3 0 s4 x2_re_a3 0 61822647521.61066
Gr2_im_4_3 0 s4 x2_im_a3 0 -56694287796.21407
Gr3_4_3 0 s4 x3_a3 0 -3849.2689865991147
Gd4_4 0 s4 p4 0 0.0034390291749299357
Fd4_4 0 s4 V4 0.17195145874649678
Gr1_4_4 0 s4 x1_a4 0 -130202809262.01865
Gr2_re_4_4 0 s4 x2_re_a4 0 -7392709157.107824
Gr2_im_4_4 0 s4 x2_im_a4 0 -29462789591.82366
Gr3_4_4 0 s4 x3_a4 0 -113591.27356952902
*
* State networks driven by port 4
Cx1_a4 x1_a4 0 1.0
Gx1_a4 0 x1_a4 p4 0 0.07071067811865475
Fx1_a4 0 x1_a4 V4 3.5355339059327378
Rp1_a4 0 x1_a4 5.282047205639696e-13
Cx2_re_a4 x2_re_a4 0 1.0
Gx2_re_a4 0 x2_re_a4 p4 0 0.1414213562373095
Fx2_re_a4 0 x2_re_a4 V4 7.0710678118654755
Rp2_re_re_a4 0 x2_re_a4 4.751370536275971e-12
Gp2_re_im_a4 0 x2_re_a4 x2_im_a4 0 2848279117741.6416
Cx2_im_a4 x2_im_a4 0 1.0
Gp2_im_re_a4 0 x2_im_a4 x2_re_a4 0 -2848279117741.6416
Rp2_im_im_a4 0 x2_im_a4 4.751370536275971e-12
Cx3_a4 x3_a4 0 1.0
Gx3_a4 0 x3_a4 p4 0 0.07071067811865475
Fx3_a4 0 x3_a4 V4 3.5355339059327378
Rp3_a4 0 x3_a4 3.5276330254138835e-10
.ENDS s_equivalent
