* EQUIVALENT CIRCUIT FOR VECTOR FITTED S-MATRIX
* Created using scikit-rf vectorFitting.py
*
.SUBCKT s_equivalent p1 p2
*
* Port network for port 1
V1 p1 s1 0
R1 s1 0 50.0
Gd1_1 0 s1 p1 0 -0.0032338265925069146
Fd1_1 0 s1 V1 -0.16169132962534574
Gr1_1_1 0 s1 x1_a1 0 -24951900993.602474
Gr2_re_1_1 0 s1 x2_re_a1 0 369935835250.25854
Gr2_im_1_1 0 s1 x2_im_a1 0 416574448141.5613
Gd1_2 0 s1 p2 0 -0.0010858199186728978
Fd1_2 0 s1 V2 -0.05429099593364489
Gr1_1_2 0 s1 x1_a2 0 27845018100.278824
Gr2_re_1_2 0 s1 x2_re_a2 0 -72943030935.58452
Gr2_im_1_2 0 s1 x2_im_a2 0 -575023015334.6757
*
* State networks driven by port 1
Cx1_a1 x1_a1 0 1.0
Gx1_a1 0 x1_a1 p1 0 0.07071067811865475
Fx1_a1 0 x1_a1 V1 3.5355339059327378
Rp1_a1 0 x1_a1 1.4471665645122728e-12
Cx2_re_a1 x2_re_a1 0 1.0
Gx2_re_a1 0 x2_re_a1 p1 0 0.1414213562373095
Fx2_re_a1 0 x2_re_a1 V1 7.0710678118654755
Rp2_re_re_a1 0 x2_re_a1 6.05836164882837e-13
Gp2_re_im_a1 0 x2_re_a1 x2_im_a1 0 1082118395574.5735
Cx2_im_a1 x2_im_a1 0 1.0
Gp2_im_re_a1 0 x2_im_a1 x2_re_a1 0 -1082118395574.5735
Rp2_im_im_a1 0 x2_im_a1 6.05836164882837e-13
*
* Port network for port 2
V2 p2 s2 0
R2 s2 0 50.0
Gd2_1 0 s2 p1 0 -0.001085819918672803
Fd2_1 0 s2 V1 -0.05429099593364015
Gr1_2_1 0 s2 x1_a1 0 27845018100.27849
Gr2_re_2_1 0 s2 x2_re_a1 0 -72943030935.58708
Gr2_im_2_1 0 s2 x2_im_a1 0 -575023015334.678
Gd2_2 0 s2 p2 0 -0.0032338265925070013
Fd2_2 0 s2 V2 -0.16169132962535007
Gr1_2_2 0 s2 x1_a2 0 -24951900993.602226
Gr2_re_2_2 0 s2 x2_re_a2 0 369935835250.261
Gr2_im_2_2 0 s2 x2_im_a2 0 416574448141.5635
*
* State networks driven by port 2
Cx1_a2 x1_a2 0 1.0
Gx1_a2 0 x1_a2 p2 0 0.07071067811865475
Fx1_a2 0 x1_a2 V2 3.5355339059327378
Rp1_a2 0 x1_a2 1.4471665645122728e-12
Cx2_re_a2 x2_re_a2 0 1.0
Gx2_re_a2 0 x2_re_a2 p2 0 0.1414213562373095
Fx2_re_a2 0 x2_re_a2 V2 7.0710678118654755
Rp2_re_re_a2 0 x2_re_a2 6.05836164882837e-13
Gp2_re_im_a2 0 x2_re_a2 x2_im_a2 0 1082118395574.5735
Cx2_im_a2 x2_im_a2 0 1.0
Gp2_im_re_a2 0 x2_im_a2 x2_re_a2 0 -1082118395574.5735
Rp2_im_im_a2 0 x2_im_a2 6.05836164882837e-13
.ENDS s_equivalent
